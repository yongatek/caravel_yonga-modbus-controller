* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_sram_1kbyte_1rw1r_32x256_8 abstract view
.subckt sky130_sram_1kbyte_1rw1r_32x256_8 din0[0] din0[1] din0[2] din0[3] din0[4]
+ din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14]
+ din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23]
+ din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] addr0[0]
+ addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr1[0] addr1[1]
+ addr1[2] addr1[3] addr1[4] addr1[5] addr1[6] addr1[7] csb0 csb1 web0 clk0 clk1 wmask0[0]
+ wmask0[1] wmask0[2] wmask0[3] dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5]
+ dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14]
+ dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22]
+ dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30]
+ dout0[31] dout1[0] dout1[1] dout1[2] dout1[3] dout1[4] dout1[5] dout1[6] dout1[7]
+ dout1[8] dout1[9] dout1[10] dout1[11] dout1[12] dout1[13] dout1[14] dout1[15] dout1[16]
+ dout1[17] dout1[18] dout1[19] dout1[20] dout1[21] dout1[22] dout1[23] dout1[24]
+ dout1[25] dout1[26] dout1[27] dout1[28] dout1[29] dout1[30] dout1[31] vccd1 vssd1
.ends

* Black-box entry subcircuit for Modbus_w_RegSpace_Controller abstract view
.subckt Modbus_w_RegSpace_Controller i_clk i_rst i_rx i_wbs_adr[0] i_wbs_adr[10] i_wbs_adr[11]
+ i_wbs_adr[12] i_wbs_adr[13] i_wbs_adr[14] i_wbs_adr[15] i_wbs_adr[16] i_wbs_adr[17]
+ i_wbs_adr[18] i_wbs_adr[19] i_wbs_adr[1] i_wbs_adr[20] i_wbs_adr[21] i_wbs_adr[22]
+ i_wbs_adr[23] i_wbs_adr[24] i_wbs_adr[25] i_wbs_adr[26] i_wbs_adr[27] i_wbs_adr[28]
+ i_wbs_adr[29] i_wbs_adr[2] i_wbs_adr[30] i_wbs_adr[31] i_wbs_adr[3] i_wbs_adr[4]
+ i_wbs_adr[5] i_wbs_adr[6] i_wbs_adr[7] i_wbs_adr[8] i_wbs_adr[9] i_wbs_cyc i_wbs_dat[0]
+ i_wbs_dat[10] i_wbs_dat[11] i_wbs_dat[12] i_wbs_dat[13] i_wbs_dat[14] i_wbs_dat[15]
+ i_wbs_dat[16] i_wbs_dat[17] i_wbs_dat[18] i_wbs_dat[19] i_wbs_dat[1] i_wbs_dat[20]
+ i_wbs_dat[21] i_wbs_dat[22] i_wbs_dat[23] i_wbs_dat[24] i_wbs_dat[25] i_wbs_dat[26]
+ i_wbs_dat[27] i_wbs_dat[28] i_wbs_dat[29] i_wbs_dat[2] i_wbs_dat[30] i_wbs_dat[31]
+ i_wbs_dat[3] i_wbs_dat[4] i_wbs_dat[5] i_wbs_dat[6] i_wbs_dat[7] i_wbs_dat[8] i_wbs_dat[9]
+ i_wbs_sel[0] i_wbs_sel[1] i_wbs_sel[2] i_wbs_sel[3] i_wbs_stb i_wbs_we o_tx o_wbs_ack
+ o_wbs_dat[0] o_wbs_dat[10] o_wbs_dat[11] o_wbs_dat[12] o_wbs_dat[13] o_wbs_dat[14]
+ o_wbs_dat[15] o_wbs_dat[16] o_wbs_dat[17] o_wbs_dat[18] o_wbs_dat[19] o_wbs_dat[1]
+ o_wbs_dat[20] o_wbs_dat[21] o_wbs_dat[22] o_wbs_dat[23] o_wbs_dat[24] o_wbs_dat[25]
+ o_wbs_dat[26] o_wbs_dat[27] o_wbs_dat[28] o_wbs_dat[29] o_wbs_dat[2] o_wbs_dat[30]
+ o_wbs_dat[31] o_wbs_dat[3] o_wbs_dat[4] o_wbs_dat[5] o_wbs_dat[6] o_wbs_dat[7] o_wbs_dat[8]
+ o_wbs_dat[9] sram_addr0[0] sram_addr0[1] sram_addr0[2] sram_addr0[3] sram_addr0[4]
+ sram_addr0[5] sram_addr0[6] sram_addr0[7] sram_addr1[0] sram_addr1[1] sram_addr1[2]
+ sram_addr1[3] sram_addr1[4] sram_addr1[5] sram_addr1[6] sram_addr1[7] sram_csb0
+ sram_csb1 sram_din0[0] sram_din0[10] sram_din0[11] sram_din0[12] sram_din0[13] sram_din0[14]
+ sram_din0[15] sram_din0[16] sram_din0[17] sram_din0[18] sram_din0[19] sram_din0[1]
+ sram_din0[20] sram_din0[21] sram_din0[22] sram_din0[23] sram_din0[24] sram_din0[25]
+ sram_din0[26] sram_din0[27] sram_din0[28] sram_din0[29] sram_din0[2] sram_din0[30]
+ sram_din0[31] sram_din0[3] sram_din0[4] sram_din0[5] sram_din0[6] sram_din0[7] sram_din0[8]
+ sram_din0[9] sram_dout0[0] sram_dout0[10] sram_dout0[11] sram_dout0[12] sram_dout0[13]
+ sram_dout0[14] sram_dout0[15] sram_dout0[16] sram_dout0[17] sram_dout0[18] sram_dout0[19]
+ sram_dout0[1] sram_dout0[20] sram_dout0[21] sram_dout0[22] sram_dout0[23] sram_dout0[24]
+ sram_dout0[25] sram_dout0[26] sram_dout0[27] sram_dout0[28] sram_dout0[29] sram_dout0[2]
+ sram_dout0[30] sram_dout0[31] sram_dout0[3] sram_dout0[4] sram_dout0[5] sram_dout0[6]
+ sram_dout0[7] sram_dout0[8] sram_dout0[9] sram_dout1[0] sram_dout1[10] sram_dout1[11]
+ sram_dout1[12] sram_dout1[13] sram_dout1[14] sram_dout1[15] sram_dout1[16] sram_dout1[17]
+ sram_dout1[18] sram_dout1[19] sram_dout1[1] sram_dout1[20] sram_dout1[21] sram_dout1[22]
+ sram_dout1[23] sram_dout1[24] sram_dout1[25] sram_dout1[26] sram_dout1[27] sram_dout1[28]
+ sram_dout1[29] sram_dout1[2] sram_dout1[30] sram_dout1[31] sram_dout1[3] sram_dout1[4]
+ sram_dout1[5] sram_dout1[6] sram_dout1[7] sram_dout1[8] sram_dout1[9] sram_web0
+ sram_wmask0[0] sram_wmask0[1] sram_wmask0[2] sram_wmask0[3] vccd1 vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101]
+ la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108]
+ la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114]
+ la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120]
+ la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69]
+ la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75]
+ la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81]
+ la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88]
+ la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94]
+ la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2
+ user_irq[0] user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2
+ wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xsram_inst sram_inst/din0[0] sram_inst/din0[1] sram_inst/din0[2] sram_inst/din0[3]
+ sram_inst/din0[4] sram_inst/din0[5] sram_inst/din0[6] sram_inst/din0[7] sram_inst/din0[8]
+ sram_inst/din0[9] sram_inst/din0[10] sram_inst/din0[11] sram_inst/din0[12] sram_inst/din0[13]
+ sram_inst/din0[14] sram_inst/din0[15] sram_inst/din0[16] sram_inst/din0[17] sram_inst/din0[18]
+ sram_inst/din0[19] sram_inst/din0[20] sram_inst/din0[21] sram_inst/din0[22] sram_inst/din0[23]
+ sram_inst/din0[24] sram_inst/din0[25] sram_inst/din0[26] sram_inst/din0[27] sram_inst/din0[28]
+ sram_inst/din0[29] sram_inst/din0[30] sram_inst/din0[31] sram_inst/addr0[0] sram_inst/addr0[1]
+ sram_inst/addr0[2] sram_inst/addr0[3] sram_inst/addr0[4] sram_inst/addr0[5] sram_inst/addr0[6]
+ sram_inst/addr0[7] sram_inst/addr1[0] sram_inst/addr1[1] sram_inst/addr1[2] sram_inst/addr1[3]
+ sram_inst/addr1[4] sram_inst/addr1[5] sram_inst/addr1[6] sram_inst/addr1[7] sram_inst/csb0
+ sram_inst/csb1 sram_inst/web0 wb_clk_i wb_clk_i sram_inst/wmask0[0] sram_inst/wmask0[1]
+ sram_inst/wmask0[2] sram_inst/wmask0[3] sram_inst/dout0[0] sram_inst/dout0[1] sram_inst/dout0[2]
+ sram_inst/dout0[3] sram_inst/dout0[4] sram_inst/dout0[5] sram_inst/dout0[6] sram_inst/dout0[7]
+ sram_inst/dout0[8] sram_inst/dout0[9] sram_inst/dout0[10] sram_inst/dout0[11] sram_inst/dout0[12]
+ sram_inst/dout0[13] sram_inst/dout0[14] sram_inst/dout0[15] sram_inst/dout0[16]
+ sram_inst/dout0[17] sram_inst/dout0[18] sram_inst/dout0[19] sram_inst/dout0[20]
+ sram_inst/dout0[21] sram_inst/dout0[22] sram_inst/dout0[23] sram_inst/dout0[24]
+ sram_inst/dout0[25] sram_inst/dout0[26] sram_inst/dout0[27] sram_inst/dout0[28]
+ sram_inst/dout0[29] sram_inst/dout0[30] sram_inst/dout0[31] sram_inst/dout1[0] sram_inst/dout1[1]
+ sram_inst/dout1[2] sram_inst/dout1[3] sram_inst/dout1[4] sram_inst/dout1[5] sram_inst/dout1[6]
+ sram_inst/dout1[7] sram_inst/dout1[8] sram_inst/dout1[9] sram_inst/dout1[10] sram_inst/dout1[11]
+ sram_inst/dout1[12] sram_inst/dout1[13] sram_inst/dout1[14] sram_inst/dout1[15]
+ sram_inst/dout1[16] sram_inst/dout1[17] sram_inst/dout1[18] sram_inst/dout1[19]
+ sram_inst/dout1[20] sram_inst/dout1[21] sram_inst/dout1[22] sram_inst/dout1[23]
+ sram_inst/dout1[24] sram_inst/dout1[25] sram_inst/dout1[26] sram_inst/dout1[27]
+ sram_inst/dout1[28] sram_inst/dout1[29] sram_inst/dout1[30] sram_inst/dout1[31]
+ vccd1 vssd1 sky130_sram_1kbyte_1rw1r_32x256_8
XModbus_w_RegSpace_Controller_inst wb_clk_i wb_rst_i io_in[9] wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
+ io_out[8] wbs_ack_o wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] sram_inst/addr0[0] sram_inst/addr0[1] sram_inst/addr0[2]
+ sram_inst/addr0[3] sram_inst/addr0[4] sram_inst/addr0[5] sram_inst/addr0[6] sram_inst/addr0[7]
+ sram_inst/addr1[0] sram_inst/addr1[1] sram_inst/addr1[2] sram_inst/addr1[3] sram_inst/addr1[4]
+ sram_inst/addr1[5] sram_inst/addr1[6] sram_inst/addr1[7] sram_inst/csb0 sram_inst/csb1
+ sram_inst/din0[0] sram_inst/din0[10] sram_inst/din0[11] sram_inst/din0[12] sram_inst/din0[13]
+ sram_inst/din0[14] sram_inst/din0[15] sram_inst/din0[16] sram_inst/din0[17] sram_inst/din0[18]
+ sram_inst/din0[19] sram_inst/din0[1] sram_inst/din0[20] sram_inst/din0[21] sram_inst/din0[22]
+ sram_inst/din0[23] sram_inst/din0[24] sram_inst/din0[25] sram_inst/din0[26] sram_inst/din0[27]
+ sram_inst/din0[28] sram_inst/din0[29] sram_inst/din0[2] sram_inst/din0[30] sram_inst/din0[31]
+ sram_inst/din0[3] sram_inst/din0[4] sram_inst/din0[5] sram_inst/din0[6] sram_inst/din0[7]
+ sram_inst/din0[8] sram_inst/din0[9] sram_inst/dout0[0] sram_inst/dout0[10] sram_inst/dout0[11]
+ sram_inst/dout0[12] sram_inst/dout0[13] sram_inst/dout0[14] sram_inst/dout0[15]
+ sram_inst/dout0[16] sram_inst/dout0[17] sram_inst/dout0[18] sram_inst/dout0[19]
+ sram_inst/dout0[1] sram_inst/dout0[20] sram_inst/dout0[21] sram_inst/dout0[22] sram_inst/dout0[23]
+ sram_inst/dout0[24] sram_inst/dout0[25] sram_inst/dout0[26] sram_inst/dout0[27]
+ sram_inst/dout0[28] sram_inst/dout0[29] sram_inst/dout0[2] sram_inst/dout0[30] sram_inst/dout0[31]
+ sram_inst/dout0[3] sram_inst/dout0[4] sram_inst/dout0[5] sram_inst/dout0[6] sram_inst/dout0[7]
+ sram_inst/dout0[8] sram_inst/dout0[9] sram_inst/dout1[0] sram_inst/dout1[10] sram_inst/dout1[11]
+ sram_inst/dout1[12] sram_inst/dout1[13] sram_inst/dout1[14] sram_inst/dout1[15]
+ sram_inst/dout1[16] sram_inst/dout1[17] sram_inst/dout1[18] sram_inst/dout1[19]
+ sram_inst/dout1[1] sram_inst/dout1[20] sram_inst/dout1[21] sram_inst/dout1[22] sram_inst/dout1[23]
+ sram_inst/dout1[24] sram_inst/dout1[25] sram_inst/dout1[26] sram_inst/dout1[27]
+ sram_inst/dout1[28] sram_inst/dout1[29] sram_inst/dout1[2] sram_inst/dout1[30] sram_inst/dout1[31]
+ sram_inst/dout1[3] sram_inst/dout1[4] sram_inst/dout1[5] sram_inst/dout1[6] sram_inst/dout1[7]
+ sram_inst/dout1[8] sram_inst/dout1[9] sram_inst/web0 sram_inst/wmask0[0] sram_inst/wmask0[1]
+ sram_inst/wmask0[2] sram_inst/wmask0[3] vccd1 vssd1 Modbus_w_RegSpace_Controller
.ends

